// System_Jtag.v

// Generated using ACDS version 13.0sp1 232 at 2021.07.28.14:45:24

`timescale 1 ps / 1 ps
module System_Jtag (
		input  wire        clk_clk,                               //                      clk.clk
		input  wire        reset_reset_n,                         //                    reset.reset_n
		input  wire [4:0]  riscv_core_0_conduit_end_disp_sel,     // riscv_core_0_conduit_end.disp_sel
		output wire [31:0] riscv_core_0_conduit_end_display,      //                         .display
		output wire [31:0] riscv_core_0_conduit_end_av_writedata  //                         .av_writedata
	);

	wire         riscv_core_0_avalon_master_waitrequest;                                        // RISCV_CORE_0_avalon_master_translator:av_waitrequest -> RISCV_CORE_0:av_waitrequest
	wire  [31:0] riscv_core_0_avalon_master_writedata;                                          // RISCV_CORE_0:av_writedata_reg -> RISCV_CORE_0_avalon_master_translator:av_writedata
	wire  [31:0] riscv_core_0_avalon_master_address;                                            // RISCV_CORE_0:av_address -> RISCV_CORE_0_avalon_master_translator:av_address
	wire         riscv_core_0_avalon_master_write;                                              // RISCV_CORE_0:av_write_n -> RISCV_CORE_0_avalon_master_translator:av_write
	wire         riscv_core_0_avalon_master_read;                                               // RISCV_CORE_0:av_read_n -> RISCV_CORE_0_avalon_master_translator:av_read
	wire  [31:0] riscv_core_0_avalon_master_readdata;                                           // RISCV_CORE_0_avalon_master_translator:av_readdata -> RISCV_CORE_0:av_readdata
	wire         riscv_core_0_avalon_master_translator_avalon_universal_master_0_waitrequest;   // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> RISCV_CORE_0_avalon_master_translator:uav_waitrequest
	wire   [2:0] riscv_core_0_avalon_master_translator_avalon_universal_master_0_burstcount;    // RISCV_CORE_0_avalon_master_translator:uav_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] riscv_core_0_avalon_master_translator_avalon_universal_master_0_writedata;     // RISCV_CORE_0_avalon_master_translator:uav_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [31:0] riscv_core_0_avalon_master_translator_avalon_universal_master_0_address;       // RISCV_CORE_0_avalon_master_translator:uav_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         riscv_core_0_avalon_master_translator_avalon_universal_master_0_lock;          // RISCV_CORE_0_avalon_master_translator:uav_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         riscv_core_0_avalon_master_translator_avalon_universal_master_0_write;         // RISCV_CORE_0_avalon_master_translator:uav_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         riscv_core_0_avalon_master_translator_avalon_universal_master_0_read;          // RISCV_CORE_0_avalon_master_translator:uav_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] riscv_core_0_avalon_master_translator_avalon_universal_master_0_readdata;      // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> RISCV_CORE_0_avalon_master_translator:uav_readdata
	wire         riscv_core_0_avalon_master_translator_avalon_universal_master_0_debugaccess;   // RISCV_CORE_0_avalon_master_translator:uav_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] riscv_core_0_avalon_master_translator_avalon_universal_master_0_byteenable;    // RISCV_CORE_0_avalon_master_translator:uav_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         riscv_core_0_avalon_master_translator_avalon_universal_master_0_readdatavalid; // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> RISCV_CORE_0_avalon_master_translator:uav_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;      // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;        // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;          // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;       // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;            // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;             // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;         // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire         rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> [RISCV_CORE_0:reset, RISCV_CORE_0_avalon_master_translator:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset]

	RV32_core #(
		.DATA_W         (32),
		.ALU_SEL_W      (4),
		.ADDR_W         (5),
		.DMEM_ADDR_W    (12),
		.INST_W         (32),
		.ADDR_W_IMEM    (12),
		.CONTROL_WORD_W (22)
	) riscv_core_0 (
		.clock            (clk_clk),                                //    clock_sink.clk
		.reset            (rst_controller_reset_out_reset),         //    reset_sink.reset
		.disp_sel         (riscv_core_0_conduit_end_disp_sel),      //   conduit_end.export
		.display          (riscv_core_0_conduit_end_display),       //              .export
		.av_writedata     (riscv_core_0_conduit_end_av_writedata),  //              .export
		.av_address       (riscv_core_0_avalon_master_address),     // avalon_master.address
		.av_readdata      (riscv_core_0_avalon_master_readdata),    //              .readdata
		.av_writedata_reg (riscv_core_0_avalon_master_writedata),   //              .writedata
		.av_write_n       (riscv_core_0_avalon_master_write),       //              .write_n
		.av_read_n        (riscv_core_0_avalon_master_read),        //              .read_n
		.av_waitrequest   (riscv_core_0_avalon_master_waitrequest)  //              .waitrequest
	);

	System_Jtag_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         ()                                                                          //               irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) riscv_core_0_avalon_master_translator (
		.clk                      (clk_clk),                                                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                     reset.reset
		.uav_address              (riscv_core_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (riscv_core_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (riscv_core_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (riscv_core_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (riscv_core_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (riscv_core_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (riscv_core_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (riscv_core_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (riscv_core_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (riscv_core_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (riscv_core_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (riscv_core_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (riscv_core_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (~riscv_core_0_avalon_master_read),                                              //                          .read
		.av_readdata              (riscv_core_0_avalon_master_readdata),                                           //                          .readdata
		.av_write                 (~riscv_core_0_avalon_master_write),                                             //                          .write
		.av_writedata             (riscv_core_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                          //               (terminated)
		.av_byteenable            (4'b1111),                                                                       //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                          //               (terminated)
		.av_begintransfer         (1'b0),                                                                          //               (terminated)
		.av_chipselect            (1'b0),                                                                          //               (terminated)
		.av_readdatavalid         (),                                                                              //               (terminated)
		.av_lock                  (1'b0),                                                                          //               (terminated)
		.av_debugaccess           (1'b0),                                                                          //               (terminated)
		.uav_clken                (),                                                                              //               (terminated)
		.av_clken                 (1'b1),                                                                          //               (terminated)
		.uav_response             (2'b00),                                                                         //               (terminated)
		.av_response              (),                                                                              //               (terminated)
		.uav_writeresponserequest (),                                                                              //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                          //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                          //               (terminated)
		.av_writeresponsevalid    ()                                                                               //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (riscv_core_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (riscv_core_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read                 (riscv_core_0_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write                (riscv_core_0_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest          (riscv_core_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (riscv_core_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (riscv_core_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata             (riscv_core_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata            (riscv_core_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock                 (riscv_core_0_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess          (riscv_core_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),          //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),            //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),             //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),         //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),        //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),      //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),       //                         .chipselect
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
